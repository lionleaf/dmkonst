library ieee;
use ieee.std_logic_1164.all;

package defs is


end package defs;
