library ieee;
use ieee.std_logic_1164.all;

package defs is

    type op_t is
        ( op_add
        , op_sub
        , op_and
        , op_or
        , op_slt
        );

end package defs;
